library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity i2c_master is
    port (
        clk   : in std_logic;
        reset : in std_logic        
    );
end i2c_master;

architecture i2c_master_arch of i2c_master is

begin
end i2c_master_arch;