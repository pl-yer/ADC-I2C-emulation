library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity rng is
    generic (
        ADDRESS : std_logic_vector(6 downto 0) := "1001101"
    );
    port (
        clk : in std_logic;
        rst : in std_logic;
        rng_data : buffer std_logic_vector(3 downto 0);
        rng_adc : out std_logic_vector(11 downto 0)
    );
end rng;

architecture arch_rng of rng is


    type t_arith_table is array (0 to 15) of std_logic_vector(3 downto 0); 
    type t_arith_table_of_tables is array (0 to 15) of t_arith_table; 
    type t_arith_mult_table is array (0 to 15, 0 to 15) of std_logic_vector(3 downto 0); 


    constant xor_gf16 : t_arith_mult_table := (
        0  => ( "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000" ),
        1  => ( "0000", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001" ),
        2  => ( "0000", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001" ),
        4  => ( "0000", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010" ),
        8  => ( "0000", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100" ),
        3  => ( "0000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000" ),
        6  => ( "0000", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011" ),
        12 => ( "0000", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110" ),
        11 => ( "0000", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100" ),
        5  => ( "0000", "0101", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011" ),
        10 => ( "0000", "1010", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101" ),
        7  => ( "0000", "0111", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010" ),
        14 => ( "0000", "1110", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111" ),
        15 => ( "0000", "1111", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110" ),
        13 => ( "0000", "1101", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111" ),
        9  => ( "0000", "1001", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101" )
    );

    constant and_gf16 : t_arith_table_of_tables := (
        0  => ( "0000", "0001", "0010", "0100", "1000", "0011", "0110", "1100", "1011", "0101", "1010", "0111", "1110", "1111", "1101", "1001"),
        1  => ( "0001", "0000", "0011", "0101", "1001", "0010", "0111", "1101", "1010", "0100", "1011", "0110", "1111", "1110", "1100", "1000"),
        2  => ( "0010", "0011", "0000", "0110", "1010", "0001", "0100", "1110", "1001", "0111", "1000", "0101", "1100", "1101", "1111", "1011"),
        4  => ( "0100", "0101", "0110", "0000", "1100", "0111", "0010", "1000", "1111", "0001", "1110", "0011", "1010", "1011", "1001", "1101"),
        8  => ( "1000", "1001", "1010", "1100", "0000", "1011", "1110", "0100", "0011", "1101", "0010", "1111", "0110", "0111", "0101", "0001"),
        3  => ( "0011", "0010", "0001", "0111", "1011", "0000", "0101", "1111", "1000", "0110", "1001", "0100", "1101", "1100", "1110", "1010"),
        6  => ( "0110", "0111", "0100", "0010", "1110", "0101", "0000", "1010", "1101", "0011", "1100", "0001", "1000", "1001", "1011", "1111"),
        12 => ( "1100", "1101", "1110", "1000", "0100", "1111", "1010", "0000", "0111", "1001", "0110", "1011", "0010", "0011", "0001", "0101"),
        11 => ( "1011", "1010", "1001", "1111", "0011", "1000", "1101", "0111", "0000", "1110", "0001", "1100", "0101", "0100", "0110", "0010"),
        5  => ( "0101", "0100", "0111", "0001", "1101", "0110", "0011", "1001", "1110", "0000", "1111", "0010", "1011", "1010", "1000", "1100"),
        10 => ( "1010", "1011", "1000", "1110", "0010", "1001", "1100", "0110", "0001", "1111", "0000", "1101", "0100", "0101", "0111", "0011"),
        7  => ( "0111", "0110", "0101", "0011", "1111", "0100", "0001", "1011", "1100", "0010", "1101", "0000", "1001", "1000", "1010", "1110"),
        14 => ( "1110", "1111", "1100", "1010", "0110", "1101", "1000", "0010", "0101", "1011", "0100", "1001", "0000", "0001", "0011", "0111"),
        15 => ( "1111", "1110", "1101", "1011", "0111", "1100", "1001", "0011", "0100", "1010", "0101", "1000", "0001", "0000", "0010", "0110"),
        13 => ( "1101", "1100", "1111", "1001", "0101", "1110", "1011", "0001", "0110", "1000", "0111", "1010", "0011", "0010", "0000", "0100"),
        9  => ( "1001", "1000", "1011", "1101", "0001", "1010", "1111", "0101", "0010", "1100", "0011", "1110", "0111", "0110", "0100", "0000")
    );

    type t_regs is array (0 to 9) of std_logic_vector(3 downto 0);

    signal regs : t_regs;

    constant x5_mult_table : t_arith_table := and_gf16(6);
    constant x0_mult_table : t_arith_table := and_gf16(1);
    
    signal nibble_ctr : unsigned(1 downto 0);

    signal rng_adc_int : std_logic_vector(11 downto 0);

begin

    process (all)
    begin
        if rising_edge(clk) then
            rng_data <= regs(0);
            if rst = '1' then
                regs <= (0 => "0100", 1 => "0110", 2 => "1001", 3 => "1010", 4 => "1111", 5 => "0000", 6 => "0101", 7 => "0110", 8 => "1001", 9 => "1010");  
            else
                for i in 0 to 8 loop
                    regs(i) <= regs(i+1);
                end loop;    
                regs(9) <= xor_gf16( to_integer(unsigned( x5_mult_table(  to_integer(unsigned( regs(5) )) ) )), to_integer(unsigned( x0_mult_table( to_integer(unsigned( regs(0) )) ) )) );
            end if;
        end if;
    end process;

    process (all)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                nibble_ctr <= "00";
            elsif nibble_ctr = "10" then
                nibble_ctr <= "00";
            else
                nibble_ctr <= nibble_ctr + "01";
            end if;
            if nibble_ctr = 0 then
                rng_adc <= rng_adc_int;
            end if;
            rng_adc_int(4*to_integer(nibble_ctr) + 3 downto 4*to_integer(nibble_ctr)) <= rng_data;
        end if;
    end process;

end arch_rng;